    localparam YES = 1'b1;
    localparam NO = 1'b0;

    localparam HIGH = 1'b1;
    localparam LOW = 1'b0;

    localparam ALWAYS = 1'b1;
    localparam NEVER = 1'b0;
